netcdf ECS {

dimensions:

model = 64, mchar = 17 ;

variables:

float ecs(model);
char model(model, mchar);

// variable attributes

ecs:long_name = "Equilibrium Climate Sensitivity" ;
ecs:standard_name = "ECS" ;
ecs:units = "K" ;
ecs:_FillValue = -999. ;

model:named_coordinate = 1 ;

:reference1_cmip3 = "Sherwood, S. C., S. Bony, J.-L. Dufresne: Spread in model climate sensitivity traced to atmospheric convective mixing, Nature, 505, 37-42, doi:10.1038/nature12829, 2014" ;
: reference2_cmip3 = "IPCC AR4, table 8.2" ;
: reference_cmip5 = "IPCC AR5" ;
: reference_cmip6 = "ESMValTool v2.0a1 (recipe_ecs.yml)" ;

data:

model = "ACCESS1-0", "ACCESS1-3", "bcc-csm1-1", "bcc-csm1-1-m", "BNU-ESM", "CanESM2",
        "CCSM4", "CESM1-BGC", "CESM1-CAM5", "CESM1-WACCM", "CMCC-CESM", "CMCC-CM",
        "CMCC-CMS", "CNRM-CM5", "CSIRO-Mk3-6-0", "FGOALS-g2", "FIO-ESM", "GFDL-CM3",
        "GFDL-ESM2G", "GFDL-ESM2M", "GISS-E2-H", "GISS-E2-R", "HadGEM2-AO",
        "HadGEM2-CC", "HadGEM2-ES", "inmcm4", "IPSL-CM5A-LR", "IPSL-CM5A-MR",
        "IPSL-CM5B-LR", "MIROC-ESM", "MIROC-ESM-CHEM", "MIROC5", "MPI-ESM-LR",
        "MPI-ESM-MR", "MRI-CGCM3", "NorESM1-M", "NorESM1-ME",
        "bccr_bcm2_0", "cccma_cgcm3_1", "cccma_cgcm3_1_t63", "cnrm_cm3",
        "csiro_mk3_0", "csiro_mk3_5", "gfdl_cm2_0", "gfdl_cm2_1", "giss_aom",
        "giss_model_e_h", "giss_model_e_r", "iap_fgoals1_0_g", "ingv_echam4",
        "inmcm3_0", "ipsl_cm4", "miroc3_2_hires", "miroc3_2_medres",
        "mpi_echam5", "mri_cgcm2_3_2a", "ncar_ccsm3_0", "ncar_pcm1",
        "ukmo_hadcm3", "ukmo_hadgem1",
        "BCC-CSM2-MR", "GISS-E2-1-G", "IPSL-CM6A-LR", "MIROC6" ;

ecs = 3.8, -999., 2.8, 2.9, 4.1, 3.7, 2.9, -999., -999., -999., -999., -999., -999., 3.3,
      4.1, -999., -999., 4, 2.4, 2.4, 2.3, 2.1, -999., -999., 4.6, 2.1, 4.1, -999., 2.6,
      4.7, -999., 2.7, 3.6, -999., 2.6, 2.8, -999.,
      -999., 3.4, 3.4, -999., 3.1, -999., 2.9, 3.4, -999., 2.7, 2.7, 2.3, -999., 2.1,
       4.4, 4.3, 4.0, 3.4, 3.2, 2.7, 2.1, 3.3, 4.4,
      3.11, 2.72, 4.55, 2.61 ;

}
